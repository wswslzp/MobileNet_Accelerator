module data_router
