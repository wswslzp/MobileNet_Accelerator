module shit #(
	parameter
) (
	input clk,
	output shit
);
endmodule
