`ifndef GNRL
`define GNRL

`define sirv_gnrl_fifo syn_fifo

`endif
